module hello_pli ();
  	 
initial begin
  $hello;
  #10 $finish;
end
  	  
endmodule
